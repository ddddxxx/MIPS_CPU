module cpu();

endmodule